BZh91AY&SY/G� ��߀Ry����ߺ����`i>�       �    P@(G�       ���  �Q�� �@�����QUc�C� oy�iT�@3��;z��  h  zzu���ޏ9�  �P ������ @F H  r���)�{�EE4 �"*��P�MiҞ"�О�=M�鐃 ��S�h
���J)?J �  #    4��d�L����L� 
���='�m&0 4   ���i�m&I�i��!����*���*1� F@2b`�z��mАVb��*���?l�Z	���;�"����
���ҥK��[G�j����r���,��%�2eK���ڶO�	P��?��)��e�QQ�B�c@
)&�%�4T�l�|��0?��iq��2�T���{1{����O��$��0�Բ�~�G���'�<�뷁�A�ID��$�$I$�H�$�"I%��D�D�H�H�$�"�I$D�����B-&��JI$�$DRI"I"H�-$I$II%�H�"I$�ZH�H��H��II$I%"I$�""�I$�$�$��D���R��������h���-�KKKD��$�$�$��D�D��D�$�IR�$�$�H�R"$��$�H�"H�"KH�"H�$�I"$��)JV����ZRZ--"I4����KE�I"Y--$����4�D�$I$�D�IRH�"$�$�$�$�"$�$�I$�$�KKJI%-$�%+JP��H�ґ$�$�$ZRI"I$��"H�I$�$�$�H�$�%)D�$�IRI$�"I$�I"H�H�"D�ZZZM-�"-&�����KK"�ih��Z"R��h���e�J$���)I$�I$�I%$�I-D�$E$�H�I$�)$�DD��DD�I�H�I"I%��D�I$�IKM)B---)4�$�I%"I""H�dI$I$I��$�H�III$DIZ$�H�I"JI$I$�$�RI"I$�$��$�%�d�%JI������ִZZM-�DZ$�H�"H�I$I$�VD�II$�ZI"$�$�KI$ID��$�H�I%�D�$I)"I-iiJR�U---&�����ZZZZD�IRI"I$�$��DMw�Yw�r��/]FV��%n�E<s,���But�(L�Hӑ�#pP��'"�M�m�����JT��Zm�Fꖓ��(�(�	c�uԹ�V[Kc)��kqԸ�jJ�m���F�ƒӋm.�[�:�X�kZ�����qĺ)�uF��T��ө�tmKm�cN�����庋�6�]i��uji��ul���Z8ғ����mն���%lun���Z�J��֥8�-Icq�[kJ����ն�:ŷ����[��q�R����qN����T��-�4�8�N��Ҥ��c�m�t���S���h�)�N:ҌKkq�$��#Jq�-*Z�ӌ[Ki.:��m�m:��Su�8�t�b�Qţ���q��mjm�)�i�N��V��)Z�YÊqE��)ũ-��SL��}ܹ��K�-֚%,q������R��iJ]6���Im���9qN�jp��K�i���8Ķ��G�cu6ێ����:���V����E�ڛu�%,m.���JKn�G�)��Iu�u�8�lm��i.��Gj:�y��%��Ɯr:�\ZT�u����u�u+Km����p�1��8u�T�-ԩ�4��%�VL%)8��c���+�����%�T��tꍺƎ��m-��luJ��4��m�h�N)��S�%��Y.���8���E8��uԺ�Ro�ƢѸ�\J��q���<�ky��R����ؗO[�:�X�[j��Kq�:�X�TҜ�R��N�R�i�4㍳�:���v�r6hѫ����rשc%F4��R�Ӎ���wb�ƚm�����4��kq�-I[�㭰�ص���:���m�V�8�KoN1�%�EDų��M�m8�;M�Ƒ�q��u�U�
1�n��8��u��N┕��n�w�J�[	��֢][g7���u&�"�7|�sw�k{kz�%Ȩ�qD����c�Lo8�Kcm�^�qM8뎥�uN�i�,����n���=uĺb�i{�8�m�\�r&5l�Ie�Q���)FZ�l��#v��^�Gb�ޛ�ӑ�8��n%�n��w3mԳ+Un���4�JT�9JK�\[M2�i%-Lm�V�8[kLum1�[q�m�-��.�t���F�K��)�,�Wih덖�jm�-)kM�[���kQn'�T����][���4ܭ����ٹqM:۶�[f�D�c9n݆�h٫r�Lɂ�̗0X(M4�\mn��eÎ1��W���I�R�4��ƱiuՒ���6�u.I��qlS�soEEG�ё��Trc���l�wM��\i�q��������H����"�O�1I���*X�Kt�������^׳�哪��8%�D�@�$�7%�=&~�z�c<���Y�Ҥ�ߋ}�ɟ*��{�Q"T���W9̨�s�������ά��R�����*9�}ܬ�G2�2�"'!UY��U���ll�seEW)\Ȋ���e��tEn9U�ݝ���Έw���މ�����U_Vw��Xʾ���VeV1�����VTDB���+2�""+2�+*�"��=��22�9�̈g8�W2��ʬ�Fg)���c�Ȫ��TOFVFer�,Fs�������D��}[��V�oV�oe�/���G2��2�2���"9�s�s)NR���̈c��U��[̪��dc��Ȏs��S��s��g+"�39NDg+2�2�ޕս��6E_f�o;�ޫ��ofVs338�+1�dG8�EUq��\�9�9U\�2��9T�s2)UJ��2�9ȆfUDVD�Uc3��s���Vg9X�s���_r�#��=������Wy�Wܾ��g9U��Ur��r����VV8�eW�#�T�ʥUr��U�Q
�c��dEW2���!�eVc�̬�*��g++9�ʩȮfDs�Dg�DeVDf|��Ϟ��Os���ޫ�ފ��3*�"Ȏs������򫏇�9ώqȆ|eVeg8Ȇs�U�Y��Vg9�;��Ȋ̥s��2!��fdDG9���XʾS3��e�os�}Y�Wܾ���z���ڻ,�F�gzdX�����s����3DD�Ffnq�Q�Ȉ�ʈ��2""��ިeUeUc*�*2�++���eeg9�T�3���W9�ܨG7�{���q�h�ު�S{7���ޞ�ob�$�*#1����fs�DD;�U��Y�Dg+��39�Q
���er"'��L��37���o2'����9̈����Q9̷�����Fg8�9��oD��̪�D�Us��w��/��ӝ��voUɔ���\ޖ/��nOh�\�黔�܍�Z�f�eW*�������y������s���|�w��[�]}w�i����#w���!�J1P�l�I��i��؈�5��G���0P��HցAl����N���5�s�[/����Ǥ�x������>>6����2&5�8��M��)Q�_)_�徬��Us���s���6��n�LK�Z�#lL��G�Ed�s܈�FUUs��Tm�1*D�m&%IJVu)�1�U9ĥ쵶�*$��T�)JII.�(�E�����!�!J�z{��܈��R�Ҕ0�J[����i%8iiLr�;	4���M���1-�)FV�D�)I)K�"Ҵ�CGJZRRcIKd��1iJԔ�fɉ0��LJ��+��B>�D��}k:Fj#�LLQ�I��TR�7�F$���ZR�/��1�%.cE�rb�ZR�4�RƢ%jTW9"�xޮDG"=�V%.�ĥ(���-)i��Z��hmiM��!KR��6���[JR��Y�%�-)GR�����6x��JN��q�TR�j��mE)�I�ĥ�����.Z&Nn4T4�Ĵ�Kf��^�JWbMS�m)n��-�E)Q�!W�R�LJR�"\��JU�1�G	JR�PJR�#��֒�L"�:�֥cIL`���M%1ؖ������2Sَ��ĥ:���q3¡\��KJ\)�X�a�%*��q�7ZS:p�R���JR�J.)�)M*�I.ќ�4p�
���e�-�)�Zc�9�	2�8��Lo��T5-)JS�C
*8�u����KCFtд�R���oP�h��9�ZLK�!��8�bVmĥ.%*�J4�)J��vKo�L�a�JPiԥ0�nq�I�d�yi�F�M����j�"�a��D��R��P�$�F���R���Zb8�Ļp�R�4l�E����JP�QIJ�LZR�uUU^�y<�s���}⒞N���i4�"vg�����^��!Ϣ"���$�"Z<$t[w���KKR�R�M�EB���I'	�Gi�d莬�Ic�qiF̊bbTT2VK�&&iIK�iJS!��1-�խk�RR��%i3��hm1.�v�b�Xѻ�1��:c�N��X��^T���XL�i{^�N=cSP��w!ל1w�'�/`蒘��A�>=<���=����s�+篑U���#�"�ވ�Ofp�W)̊�g9�Gz�����z��Ug1�3�dG1���O;ʬ�g1UY�TUs��Cy=̞��9��1\q�s=���w{{9���r��r�=���ފ��V�y|�ew�Q1��ȅg��LVDDc��r��{1�ʩ��r��c�z��7�����:���ĝ���5�۠���G�a�.0�� �o462Z0���FH�Idđ��5���}�a1B��R.�$�ě���E�?#�4�)��-+S#��z�#�Jȍ�Ȋ�⸎B�{y��0F8�Q��C�����aVx�p�RT.>>���ԛ��t���EE&N4|`�g�ȏ�:a���TT$��c�%F��w/-�'-��I��L/�:t�	���l���~0�mN?<l��i̍�e,��"�x��0�b���Q�aDY[.!H���d�Ŧ�1�Sʍ��G��O�$��fEa��?8��*#Ȫ��OEDoz�1�����q�1��ϱ��Ǝ�l�\"O�:zl�l�c㥘LL6~�"<���~�d��K�=�wIu�c~=�F���]���0���zLF����(S��m-�ҏj�
,�������g�l�'d��E���ĸ�oO6�n'f�m�(٢c�!Ç�	��Y͜�ކ�,�PY#�~q����m��M�ۘ�mM�%�GL�K��S!�0�B���c��Qޥ7�2��5�F�S���6a�a����h����)C.c�����C�?[�4�8�3��_#ф�4'�*#
?�$����.���Chot1x��0~���Վ�N���Ɩ�"�i�)�?�4�Qn8����i�<�����6�6�\R�c�4��<�T�Vۭ�R��Ĵ��[y-��ͻ�DZx�
i��4ߙ��m�4�-�&...��er�q����Ǟ�4�1�6���n��ߣ"cQ��|��,�������$������udՂhn��8n�dn�&�hw��e���[:ȒM�:I�Z�dѪ��m:4�n�23��F֧+I��w�j��kL2NS!�	$F�6t���a�e][��sG3*na��H�H�K<ۄ��I5�+L8�p���f�d0�r���ht,M�FCcsU|L.5	��Th��p��|dyn�k�Q��1���ڔ�ª>���G9
��B��R�#yL�22;�M�{\0�#	��j ���9�Y�t:��9�s���$��fJ"�2>��0�0�i�Ȋ#�NB�ѷ���|ӎQ��	q���* ���'ċ$}	8Ibb$�K&Q�u7�����9C���h�D��:�#"��6۵�y���q2t1:�8�62�9���չ�0���2�fM��橹����9�)�v>(�$�H�ϛq�4�i���X5w1hm2�\gy���"f6�HȑD�0�`ِ�0�qh5�L��	6�q��cqG������Q���W"7���)�9H�o/�����z"�gzd��/�c{zc���>��Sj`po5�%��jl27�hˑ���S��r4v;�s'��t,N�֧I�ww6���R��)���~���dD~��CGaD͍&�N�CUr��cB��AC�p��~0�N�E�">�I��2(�Q��~�i�����Z�q����:I��r$zl���FBN,�<x�pEt��J��q!H{��q3O�-o�������uk:�q�K�������P��h����FQ&�p�AD~$�$��l��D�"E�O���I��D`n��� -�$;.T�;�ݥ�؊�)�6�d���y��Imou,bR�V�o�m�3�R�mo).:�T�%ǜJZK�%�b]u���4��SʊSM4K�'o3�*ۖ�8��{��).&���{y�)F�iO���R\�ƢT�%ǜJZK�&<�o�-�j��R"�KQ��E�!��|�7Vry���?	����UVV9�Ȩ�r'���}��R""���ʈ�DTs*�\��{3��eF9��defFV;ѽ}��DW3#�YY�U�c""�����Fc9�V"+��W2#��ޮ����}\�U#�\̬����W{!Y��TUr9�Q�}|�f���"���S����{��͛����ie�P�� }A�l�8�	`(v�h���h�;�;�F�x0�0�Js�W6T�š�J�b9�Yao��p�sm��W1w�����Ȉc2'�LoR������_;��?�sq��F�2������I�xa�qZ-�7���%���j$���>�$�r$��D�Ɲ���M6�.6�l�����w�U�����Y`�1$�,J2"��Du�O�K��k&�	���b����9Z��D�%����N21h�~���&=�Ě.�
'�h��~0�ND��8~><j:N���y�8�X����q��=B!��G��H�F���7��,�,�O��m0���ݶ��qIQ)J��0��0������VDe'����11)�T\dxB�Y�FLG����0��:u1��2�æ�>��_��Z͊4\.U�hP�
�4�����6H���Z&~<p��L&9Q�%B%�aƟ1�1�}�4���gG"8�DCG�."��J�t�h�\|IE�>~Z[i�6���X��	D��O���O�2��c���r0�|ll���F�U�}e���R���ȥ�S!�#��r#���*�7����!��T��s��<�>�MS#Sc����fε�,��b����
,����ц�ÇV���)i�-M1ڷLd�&'6SJ�S��А��0�dĖY����F���p�GM�dl�h�fe��<�"�4���T��GYR�4�bT�M��Z�m�,��[�<��㍺�c�إ��n��i.%k>~m�m��Lm)i��u�q�)֭.��q�V�TiN���-1�����q8ښ��c�u��jx���W#��J�m�8�����a���X�$j`��P�a4�pJ�&իU�ǅ����V�v\0t$�DDh�#"����Fa�U����pl��?G��	E��}�P�>(���[O�<���|�M:�wln&:uƚ~�va3PÁg���	0�P�E�g!�!��������M4�#�W՝쌌�����g#�}L�2�#���Ee_orX�����1���y�����%�0��C ��Cő�A�����Ƣ�a�"!��f9���6�ͩ����q-9*��-�7Aq$h��2Q�E�,���??C!��Ӂ��˂��S����U�JK�gN�$��(����g�L�C�T$},�6~�!�b" h���o��mǶ[q�%�У��QQӰ���8|~:x�v<Nˈ|j&J���Ψ��y8���^E5/����W[�1,)L�QeF�3��g";���\VN$��d2-���h�F�����C�*|TD\E��$��}�0�a�������6��TK�9�Ը⸕���>>2&>?h�=
<}LEÄ����:l���柖�6���m����������E��8va(�Gv��c�Y*~y���7����i�7DGa�B�r��.Gc{y�:���O�\L$�~��8��Q�ϟ�㭱�i~)��oƔ�ͥ�Zuؔ���S�m��4�.��K~q�b�moѷ��4�O��i��z(��/:��Jm����=io�%�����Jy�#�uȗ��n�S�m���W�i*y/��bJy������f�_��ͼ�Zy��Q�]I�ιk�>����y%))d�
ZV�e�*;���ʱ��G;��̮dUr1�Q�r��O_;��Vz9U\��C**9����_w�s)FeS#U�es���b{�H��ER����㜊�yW�FEVdg8�C29�r3�}ʫ���3UG9��Z��9��9��7��I#+��\��W'�}��H��Wܞ�Һ�OZɑ}���o�=s���C�G�dxp��7�$n��4�d�I��i$�$�����G�k,"Ŗ���e�L�f�GI���H��r��{�,�R�S!��D!��8�b�Qʥ9�討to"Wo_}�A�!���&#Q�0�:P�����%}g	�#f��0�Ȓa�゜K��%N���A��&�Bc!����Ϗ���8hr9
D�E�~??8��N8��8�8���7Cp�$Ӏ�M�[$p�n�\%���P�P�&��[�?$�1lr�H��?�
>�;���7��s�����kW����xC�.Bߟ��D�ԕ�ݟ�K�����2�XZI0ޥ1�Q�UDS{���1RfBVIp��G�$DF�6bE���m.219�'Se�
Y���L4n:��#Kkuӎ)��\m�N����Q�|L?4j"�8^�GNG���%G��a��N>[y�8�q�8���$��a�~?C��C�K�-��J˅%ڋ��)	ȳ
&�?a"MG�E��,��E�ҡ������kZ�1��J_�TF;�fDoUFTo8�"��q���q��e7�{*�؈�Q
�5�d'	;���#���|L([�&:}�0�g��+M��?4��m��T.9�8��~TQ$�BĒY��".&" $�������cP�$�?C�:?E#��eT��|�O������S�~b�[�~x��\<ǜTy�K��<����^R��^J�둎6�T�w�o(����FDJ�{F�^4ל��_a�n��sP�N�َ�G�u�X��mǔ��v<ړoK�b]o�Em.�$�i�K9'k";c�,�G{psv���ъe�Ma9�vƛ2�D�bZ�2e���ϡ�s��޹͝0șaP��l�heӸF2`ɱr����n�D������zl��x�D�D�p�_va�Ȋp��y��[��1�o��m�v:���JZڅ0��ʊ��rg�To+ѽ�V���N���oEN����8ee��͍	̕h�iNf����[���u0�OC��D�ǝb\R�i��-']qQ���v�������|t�0�D&0�l�2"�8|���tǘ�o�)Ƣc�q�]q���I�J�Z<p�0�c�9$�e��aP٨�mN��[#գQ���fG���?Bf0���-��Q~?0��l��q��%I_Δ�&\l��%�ݖ�ȓ�IKS"9�̈�!�ޥ1�Jcz��r�)������b0�Y���(��0�R|T:Y��ό��9�0�m�ߖҒ�R�������i���ߴQ��t�_F�:a��çA��am�F<�+��q2�~.;a���p��F"K,��t��(��dEu.4��\-�L~qm6�U�\�1ƴ�㑆ύ�4Q�ş��-�¡'J,�&a2�ߞ~b�i��>cM�����cKN�/፸y.�N��αo(�J�<�JKuKt�ιiSӏ24Υ�:�lN*<im4��ZX��ĽIK;�q*��Ǖ�G-r�N�\m��j�YSy�c����Nڗi���>UDr9̧+9Yʎl�fO[����odeEB#��C�s�ʪ���OOV����r�W+��U�R�y��feg2����s��'�����fOTDq��9YY�VW33�s3����G�g#ѓ��"��̮�9[׽}�9�s��UG9Q���{��}�;�VDo29Q��򢙙S��Er��}��]}̞��Ȟ�7�7�k=�G�Oz{�O>�� �%=`�c\Q:���L7������b�TK�1�K!�%f8�G;����VD�f7�c�/�f�0цC?C}$�F>�*�.	0�>>���Q�KG_�K��[���-Kq�J�CE��F�F��z&Y0�4|a�0�Q�L|h�٨�����mǛm�Ҕoq��i1�j���Kx��8~0�a�g���$՟����\y/�m�\r<����W��0�gc	��}	>>.#�:l�|h�r"�G�Q>R_8�<��lJ���F�9���Xd-��Y�!Q�w��FTw��Tv�����^���q��'�o{�q�f�)�
��	t����FΙ	�7Z^J����%�i�5�<n:|d.,~-~�O�������Bcȋ�Ӭ-������!�&�����ٳ����I0�>�p�Q��u����0�ZkM��=.F?<��	9�$����a�9B������E�T.>m�w�Ck|��Ɯi-)q)Z��1e�0�̄8���)=LUR�����50ц���~�Ѹh�\>�����Q#P���!�p��?d%�ǡ�����R?8��Թ8�FG8��:�СOC
.鐣�Cg�##B��H�%孊m��|٧�j#m�oͼ��:�p��ic���ږ�Rq-?1���q�K��m��Sf)�c��iKZV�<m��1�%�u�[4�7�-��i�c�?^�y��Im��\R܉K�i�?7
��#~�N�i��h�6�4��i�j.5S��qM�\i/�N��Ǡ�%���B]���1�3�.t��v�:l�z#	�a�p���Dn�T&(�^4��S�M�i�n.0������|a��$�h��1�̎o�0�`��P��KJq�_�;��oT�V��)*��Ȏ7�̈��G�G�U#y=
aK�%g{{��{��T�\*�K��Q4�		IHK����A�Tj��.Ř2�	u��x�n8�8��������*2x�Yu����x�!8I�p���zLl���?>y��u�ɭ���lA��ۑ�!n�*��ht��5�<Vp�ό�y/,���ȵŽ��a�bMC�ç���b8x��f~(�,�M�R*0ŭ��aS>���(�y\Ȋ�c���g��c�Eoz�V�۽�qfd'	��!GOŰ��3�ř��������Bb8p���s[E�li,�di�O>?C	��*L���o�&�Z-�R��iL�a�������ߋ�G�N�2���aӥl�F%Զ�V��4����ǡ�ӆ�&���Ŝ,��	�TB�E��:�?:�柍��ZQU�u�iƛh�OuO�jJR�o8����qן�m�m��⎴���h��q.<�~���<ڊR��z1���6Ѹ�_�K�����%�ǜTp���屦���r$�_jUy�1E*)�Ns'���T�켈���Vg"��Q�G8��R��"8�o7�U��s�������3���;�+"��Ȭ�2\�s�]�辞�oW+"�����+��V*yY��r9��s"Ȏs�3���o9�]�U^w���39YȬc/�Q=����fTr�+8��B���'����k��{���� ��Zգ+%�6�U�n�t��Sr6r6K��Z��	B�	��D�����z9�U_=��Vw��ʍ�dG�q��q�odLc�_dD�ow���<�b���� ���a�0�Y(z>?����C�>�����+\TZ_�&$٣��6z<t��b,���0���G�z_~}�|�)�K�>�K����0م<�h���?LGK8Q�cŔ~L'Q�͑�>6t�D����_��0��h�g�\4aGOŌ?4��?6���Ӱ민�]u������VE(��(�j%��DS���R�#Њw�W�3��8�by�S�S�&BJ�Y'�?|���C!��;4�R��Z�jRJ}���,�I$Y'����0�?)H������ZZ\i�-�����D���O�	,�����=�ce�#�aG孷��-���7\?G��d�G�G��?C%7M��
��>(�,m.����Қ{m���R�[��g+;�\�2'��ST�w)��;�L����̆4dd0�|p�TCFY��g!��7?Fp�G��m>[6��%�6�M��i�t����m�ّ��h�4~8~�K������LlȶߛiJz6��y�Z�|�%&�SKc�p�8�Kv���ji+d��]i���i�~Ko-ƞc�><����4�֤��/�<ǟ���R�SK�c��:�?:�uK[��&7�6���-֖��.Gb����}�%|y�b[EƢ��~�~[���~���??4i��KRR�c�z<ǟ�=�uM-�����&Y2j��磶�i�m�Sc��M1�C�v�7��\�"��I)&$�S���:�8cMj�1��XML2q2�I����r�5L���\��F�h�0�$ѐ��ξKLmlK�h~B`T�<v5�8|zH�l|T;
$��#��d��IDn%��1�2;�Ur��VT8�Or����9Q[�S�Do2�����Sw��������DU{ʌ��Ȭ`\qqhѱ�����&�^���,�p��	�2}I'���#lr-�GSjJR�Li��iIJZC��m0!����2�
�0�E?C	��r��FʆB��KM����2I��� �%|t��6d#��ӱ�Bp�z���c��E�.�Xp٦�u��TW&J��nh�:/"[j�0��.*����
4��|�Ҵ��G������q��+[Ц9ʮ9�Sz��w��toD�oou���Jq�A�>��K'���0�T6I��	Y��#G�rd'	(�>?��-�6�NV�ߒ��Wj���_�G����$dä�Ο�C��t�GJ,�����)�S6q%��8|~0�b$��QD�Ȋ��î���:��1,�i���V�昖BZ�}�I?��G#gC���h�R?��O�]̝vv�[�>a�i��/���1��9���UUT��d�lͱ���{�TG�?B�}Q�EIl��dk5J$��#�O�(X�H/�"�lk��NL�c]��-�ي�I1�&0T�6P�b�c'�v�8�f����b�Yd&K�ڪ$ݮZ�9�!U�SVT���*7oƶ�q�Y��G\A�lhI��%r��ͅ��i�u�[ϻ��vZ(�-�U��PKK�؃����!R��@��I,��H	��Q)�#��O�W�3�;� �=�C��i��N_����р{!<Cd���K$�sD��_����_�o&��I�'1<i����m:�O-�m��9�c��
�d���w|��T~L~K��OB����~s��4*�ХR��zd�Cb��ܼ�����&[��r�蟹7�Y=��3��_O������6v�N��>�|�.�L'����`����I������2��&��쾹��]�)��r�㓼�ss�����-<2٨n���&�����ɩ��_�3��E��Q.�	nV��v�aHL������q�"��04O	B$��|�i'9�H�"����$jljf[l�I����#i��9L�aB��Մ�2�-��m�cl��[nh֍�-�l�֋"ȴF�-�b,��F�k[i��4M�F�E�k�Y��Y,��F��n�[b����6fE���kZڋBdY��3dM�-�h�l���d"-�֊,�[�d(�-mE���E���k�d�Kl�VQ-��"дMF���DE�mF1&ֶe�m���ׅ����Z%%(��s����q��%W���̕�ʤ��E�B�]����b񹉁�d�P���}bȦ�ޝɭ+a�/?�bwm)���x^�Z���A7*��{	>$Oz�y��v�Mҁ
�AN
Q}T����qO6;��_��/~��l�r`��L�~������%��:E�O�_���O��z_9���Y8W��.��=i��O9����R���5��S�;�Q���a`X �c�=�4�O�w�0<R�*���$}���`Ną;ǜ *�������|_�X^f?*̯��1{$K)�PI�b�i	��0��z_�ί�z�
�sNs�}̍�x��&ɩ���N*�<_{7C�����oSv.�&�V�+�i40���X���/�i8�qqb�5V��u����5��o>���f�L':9�T�������������uY��r�Z{�*^��9�_dv?:N��)~'�w��g��7Ngy ?����vN��yq���/�<��:Y�՘�֧�^��훯�z��d�{RQ󎞏xݺU����&���ķ��Z���ا�|!*ZC�ܜO|ɧ����su��>s��W�j.C�x8�)���&8X|���i3�Y��ΛL�,��O���ybxO�u�<o�O���V��[ j@�a�J	)jh��М��l��Zd���W�x���T%K������Le��2zM���L���qmOE��W"���m�Mש��N) \n/W��{f�œ�ޜר�ΓS�<I�s��:���N�v�{�reER�L'��}���.�ܝ���&O��꾏	��6MWGj�������IS���T��&w��>�:����s}r���WW���<���"�I�\�_�>dN�]��B@�